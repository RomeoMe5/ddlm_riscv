module top (SW, KEY, LEDR);

    input wire [9:0] SW;        // DE-series switches
    input wire [3:0] KEY;       // DE-series pushbuttons

    output wire [9:0] LEDR;     // DE-series LEDs   

    b9_6bit_dec_mips_maindec dut (SW,LEDR[0],LEDR[1],LEDR[2],
										LEDR[3],LEDR[4],LEDR[5],LEDR[6],{LEDR[7],LEDR[8]});
 
endmodule

